//      // verilator_coverage annotation
        //========================================================================
        // Integer Multiplier Simple Implementation
        //========================================================================
        
        `ifndef LAB1_IMUL_INT_MUL_SIMPLE_V
        `define LAB1_IMUL_INT_MUL_SIMPLE_V
        
        `include "vc/trace.v"
        `include "vc/counters.v"
        `include "vc/muxes.v"
        `include "vc/regs.v"
        `include "vc/arithmetic.v"
        
        module lab1_imul_IntMulSimple
        (
 069399   input clk,
 000001   input reset,
 007090   input  logic        istream_val,
 007090   output logic        istream_rdy,
 000293   input  logic [63:0] istream_msg,
        
 007090   output logic        ostream_val,
 007083   input  logic        ostream_rdy,
 000771   output logic [31:0] ostream_msg
        );
        
 000293   logic [31:0] a;
 000759   logic [31:0] b;
 007090   logic        next_ostream_val;
 000771   logic [31:0] next_ostream_msg;
        
          assign  a = istream_msg[63:32];
          assign  b = istream_msg[31:0];
        
 034699     always_ff @(posedge clk) begin
 034699         istream_rdy <=1;
 003545         if( next_ostream_val )begin
 003545           istream_rdy <=0;
                end
               
 034699         ostream_val <=next_ostream_val;
 034699         ostream_msg <=next_ostream_msg;
                
            end
            
%000000     always_comb begin
%000000       next_ostream_val = ostream_val;
%000000       next_ostream_msg= ostream_msg;
 007090       if(istream_val && istream_rdy)begin 
 007090         next_ostream_msg = a*b; 
 007090         next_ostream_val = 1;
              end
 007102       if(ostream_val && ostream_rdy) begin
 007102             next_ostream_val =0;
              end
            end
        
        
          //----------------------------------------------------------------------
          // Line Tracing
          //----------------------------------------------------------------------
        
          `undef SYNTHESIS
          `ifndef SYNTHESIS
        
          logic [`VC_TRACE_NBITS-1:0] str;
          `VC_TRACE_BEGIN
          begin
        
            
            $sformat( str, "%x", istream_msg );
            vc_trace.append_val_rdy_str( trace_str, istream_val, istream_rdy, str );
        
            vc_trace.append_str( trace_str, "(" );
        
            $sformat( str, "%x", a );
            vc_trace.append_str( trace_str, str );
            vc_trace.append_str( trace_str, " " );
        
            $sformat( str, "%x", b );
            vc_trace.append_str( trace_str, str );
            vc_trace.append_str( trace_str, " " );
        
            $sformat( str, "%x", ostream_val );
            vc_trace.append_str( trace_str, str );
            vc_trace.append_str( trace_str, " " );
        
            vc_trace.append_str( trace_str, ")" );
            $sformat( str, "%x", ostream_msg );
            vc_trace.append_val_rdy_str( trace_str, ostream_val, ostream_rdy, str );
            
        
             end
            `VC_TRACE_END
          `endif /* SYNTHESIS */
        endmodule
        `endif /* LAB1_IMUL_INT_MUL_SIMPLE_V */
        
