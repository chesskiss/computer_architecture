module hello;

initial begin
  $display ("Hello");
end

endmodule
